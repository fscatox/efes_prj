/**
 * File          : tb_ps2_controller_pkg.sv
 * Author        : Fabio Scatozza <s315216@studenti.polito.it>
 * Date          : 29.11.2024
 */

interface ps2_if;
  tri1 clk, dat;
  bit clk_od, dat_od;

  // device drivers
  assign clk = clk_od ? 'z : '0;
  assign dat = dat_od ? 'z : '0;

  modport dev (
    input clk, dat,
    output clk_od, dat_od
  );

endinterface

package tb_ps2_controller_pkg;

  timeunit 1ns;
  timeprecision 1ns;

  //
  // Randomization utilities
  //

  function automatic int unsigned lfsr();
    // any non-zero seed
    static bit [31:0] state = 32'hAE1F_B42C;

    // XNOR Taps: 32,22,2,1
    // https://docs.amd.com/v/u/en-US/xapp052
    state = {state[30:0], ~^{state[31],state[21],state[1],state[0]}};
    log("LFSR", $sformatf("state = %0d", state));

    return state;
  endfunction

  function automatic int unsigned lfsr_range(int unsigned maxval, int unsigned minval = 0);
    return minval + (lfsr() % (maxval-minval+1));
  endfunction

  //
  // Logging utilities
  //

  function automatic void log(string who, string what);
    $display("[%0t] [%s] %s", $time, who, what);
  endfunction

  function automatic string flagsToStr(ps2_pkg::flags_t flags);
    unique case (1'b1)
      flags.frame_error: return "frame error";
      flags.parity_error: return "parity error";
      flags.clk_timeout: return "clock timeout";
      flags.rqst_timeout: return "request-to-send timeout";
    endcase
  endfunction

  //
  // Device model
  // See: IBM PS/2 Reference Manuals, Keyboard/Auxiliary Device Controller, 1990
  //

  class Ps2Device;

    const time tclk;
    const time ts; // from data transition to falling edge
    const time dt; // clock shift

    typedef bit [7:0] payload_t;

    virtual ps2_if.dev ps2;
    bit clk;

    function new(virtual ps2_if.dev _ps2, time _dt = 0);
      tclk = 50us;
      ts = lfsr_range(25,5)*1us;
      dt = _dt;

      ps2 = _ps2;
      clk = '0;
    endfunction

    task run();
      ps2.dat_od = '1;
      ps2.clk_od = '1;

      fork

        begin : clk_p
          #dt;
          forever #(tclk/2) clk <= ~clk;
        end

        forever begin
          @(posedge clk);
          log("Ps2Device", "Checking the bus state");

          if (ps2.clk) // not inhibited
            if (ps2.dat) // not a request-to-send
              _tx();
            else
              _rx();
        end

      join
    endtask

    task _tx();
      payload_t py = payload_t'(lfsr_range(2**8-1));

      bit [10:0] pkt = {
        1'b0, // start bit
        {<<{py}}, // payload lsb-first
        ~^py, // odd-parity
        1'b1 // stop bit
      };

      log("Ps2Device", $sformatf("Sending '0b%b' as '0b%b'", py, pkt));
      foreach (pkt[i]) begin

        // Generate bit 't1' before the falling edge
        #(tclk/2-ts);
        ps2.dat_od <= pkt[i];
        log("Ps2Device", $sformatf("(i = %0d) ps2_dat <= %b", i, pkt[i]));

        // Check for inhibit at every falling edge, before generating
        // a transition on the bus
        @(negedge clk);
        if (!ps2.clk) begin
          log("Ps2Device", "Clock collision: aborting tx");
          ps2.dat_od <= '1;
          return;
        end

        // Generate the falling edge
        ps2.clk_od <= '0;

        // Generate the rising edge
        @(posedge clk);
        ps2.clk_od <= '1;

      end
    endtask

    task _rx();
      payload_t py;

      for (int i = 0; i < 11; i++) begin

        // Move to the sampling point
        #(tclk/4);

        if (i > 0 & i < 9) // data bit
          py[i-1] = ps2.dat;
        else if (i == 9 & ps2.dat != ~^py) begin
          log("Ps2Device", "Host parity error");
          $stop;
        end
        else if (i == 10 & !ps2.dat) begin
          log("Ps2Device", "Host frame error");
          $stop;
        end

        // Reverse roles for generating the acknowledgement
        if (i == 10) begin
          ps2.dat_od <= '0;
        end

        // Generate the falling edge
        @(negedge clk);
        ps2.clk_od <= '0;

        // Generate the rising edge
        @(posedge clk);
        ps2.clk_od <= '1;

      end

      // Revert acknowledgement
      ps2.dat_od <= '1;
      log("Ps2Device", $sformatf("Rx done: '0b%b'", py));
    endtask

  endclass

endpackage
